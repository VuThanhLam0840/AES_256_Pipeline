module sbox(
    input  wire [7:0]  index,      // Input byte (0-255)
    output wire [7:0]  out    // S-Box output
);

    wire [7:0] sbox_data [0:255];
    
    // S-Box lookup table
    assign sbox_data[0]   = 8'h63;
    assign sbox_data[1]   = 8'h7c;
    assign sbox_data[2]   = 8'h77;
    assign sbox_data[3]   = 8'h7b;
    assign sbox_data[4]   = 8'hf2;
    assign sbox_data[5]   = 8'h6b;
    assign sbox_data[6]   = 8'h6f;
    assign sbox_data[7]   = 8'hc5;
    assign sbox_data[8]   = 8'h30;
    assign sbox_data[9]   = 8'h01;
    assign sbox_data[10]  = 8'h67;
    assign sbox_data[11]  = 8'h2b;
    assign sbox_data[12]  = 8'hfe;
    assign sbox_data[13]  = 8'hd7;
    assign sbox_data[14]  = 8'hab;
    assign sbox_data[15]  = 8'h76;
    assign sbox_data[16]  = 8'hca;
    assign sbox_data[17]  = 8'h82;
    assign sbox_data[18]  = 8'hc9;
    assign sbox_data[19]  = 8'h7d;
    assign sbox_data[20]  = 8'hfa;
    assign sbox_data[21]  = 8'h59;
    assign sbox_data[22]  = 8'h47;
    assign sbox_data[23]  = 8'hf0;
    assign sbox_data[24]  = 8'had;
    assign sbox_data[25]  = 8'hd4;
    assign sbox_data[26]  = 8'ha2;
    assign sbox_data[27]  = 8'haf;
    assign sbox_data[28]  = 8'h9c;
    assign sbox_data[29]  = 8'ha4;
    assign sbox_data[30]  = 8'h72;
    assign sbox_data[31]  = 8'hc0;
    assign sbox_data[32]  = 8'hb7;
    assign sbox_data[33]  = 8'hfd;
    assign sbox_data[34]  = 8'h93;
    assign sbox_data[35]  = 8'h26;
    assign sbox_data[36]  = 8'h36;
    assign sbox_data[37]  = 8'h3f;
    assign sbox_data[38]  = 8'hf7;
    assign sbox_data[39]  = 8'hcc;
    assign sbox_data[40]  = 8'h34;
    assign sbox_data[41]  = 8'ha5;
    assign sbox_data[42]  = 8'he5;
    assign sbox_data[43]  = 8'hf1;
    assign sbox_data[44]  = 8'h71;
    assign sbox_data[45]  = 8'hd8;
    assign sbox_data[46]  = 8'h31;
    assign sbox_data[47]  = 8'h15;
    assign sbox_data[48]  = 8'h04;
    assign sbox_data[49]  = 8'hc7;
    assign sbox_data[50]  = 8'h23;
    assign sbox_data[51]  = 8'hc3;
    assign sbox_data[52]  = 8'h18;
    assign sbox_data[53]  = 8'h96;
    assign sbox_data[54]  = 8'h05;
    assign sbox_data[55]  = 8'h9a;
    assign sbox_data[56]  = 8'h07;
    assign sbox_data[57]  = 8'h12;
    assign sbox_data[58]  = 8'h80;
    assign sbox_data[59]  = 8'he2;
    assign sbox_data[60]  = 8'heb;
    assign sbox_data[61]  = 8'h27;
    assign sbox_data[62]  = 8'hb2;
    assign sbox_data[63]  = 8'h75;
    assign sbox_data[64]  = 8'h09;
    assign sbox_data[65]  = 8'h83;
    assign sbox_data[66]  = 8'h2c;
    assign sbox_data[67]  = 8'h1a;
    assign sbox_data[68]  = 8'h1b;
    assign sbox_data[69]  = 8'h6e;
    assign sbox_data[70]  = 8'h5a;
    assign sbox_data[71]  = 8'ha0;
    assign sbox_data[72]  = 8'h52;
    assign sbox_data[73]  = 8'h3b;
    assign sbox_data[74]  = 8'hd6;
    assign sbox_data[75]  = 8'hb3;
    assign sbox_data[76]  = 8'h29;
    assign sbox_data[77]  = 8'he3;
    assign sbox_data[78]  = 8'h2f;
    assign sbox_data[79]  = 8'h84;
    assign sbox_data[80]  = 8'h53;
    assign sbox_data[81]  = 8'hd1;
    assign sbox_data[82]  = 8'h00;
    assign sbox_data[83]  = 8'hed;
    assign sbox_data[84]  = 8'h20;
    assign sbox_data[85]  = 8'hfc;
    assign sbox_data[86]  = 8'hb1;
    assign sbox_data[87]  = 8'h5b;
    assign sbox_data[88]  = 8'h6a;
    assign sbox_data[89]  = 8'hcb;
    assign sbox_data[90]  = 8'hbe;
    assign sbox_data[91]  = 8'h39;
    assign sbox_data[92]  = 8'h4a;
    assign sbox_data[93]  = 8'h4c;
    assign sbox_data[94]  = 8'h58;
    assign sbox_data[95]  = 8'hcf;
    assign sbox_data[96]  = 8'hd0;
    assign sbox_data[97]  = 8'hef;
    assign sbox_data[98]  = 8'haa;
    assign sbox_data[99]  = 8'hfb;
    assign sbox_data[100] = 8'h43;
    assign sbox_data[101] = 8'h4d;
    assign sbox_data[102] = 8'h33;
    assign sbox_data[103] = 8'h85;
    assign sbox_data[104] = 8'h45;
    assign sbox_data[105] = 8'hf9;
    assign sbox_data[106] = 8'h02;
    assign sbox_data[107] = 8'h7f;
    assign sbox_data[108] = 8'h50;
    assign sbox_data[109] = 8'h3c;
    assign sbox_data[110] = 8'h9f;
    assign sbox_data[111] = 8'ha8;
    assign sbox_data[112] = 8'h51;
    assign sbox_data[113] = 8'ha3;
    assign sbox_data[114] = 8'h40;
    assign sbox_data[115] = 8'h8f;
    assign sbox_data[116] = 8'h92;
    assign sbox_data[117] = 8'h9d;
    assign sbox_data[118] = 8'h38;
    assign sbox_data[119] = 8'hf5;
    assign sbox_data[120] = 8'hbc;
    assign sbox_data[121] = 8'hb6;
    assign sbox_data[122] = 8'hda;
    assign sbox_data[123] = 8'h21;
    assign sbox_data[124] = 8'h10;
    assign sbox_data[125] = 8'hff;
    assign sbox_data[126] = 8'hf3;
    assign sbox_data[127] = 8'hd2;
    assign sbox_data[128] = 8'hcd;
    assign sbox_data[129] = 8'h0c;
    assign sbox_data[130] = 8'h13;
    assign sbox_data[131] = 8'hec;
    assign sbox_data[132] = 8'h5f;
    assign sbox_data[133] = 8'h97;
    assign sbox_data[134] = 8'h44;
    assign sbox_data[135] = 8'h17;
    assign sbox_data[136] = 8'hc4;
    assign sbox_data[137] = 8'ha7;
    assign sbox_data[138] = 8'h7e;
    assign sbox_data[139] = 8'h3d;
    assign sbox_data[140] = 8'h64;
    assign sbox_data[141] = 8'h5d;
    assign sbox_data[142] = 8'h19;
    assign sbox_data[143] = 8'h73;
    assign sbox_data[144] = 8'h60;
    assign sbox_data[145] = 8'h81;
    assign sbox_data[146] = 8'h4f;
    assign sbox_data[147] = 8'hdc;
    assign sbox_data[148] = 8'h22;
    assign sbox_data[149] = 8'h2a;
    assign sbox_data[150] = 8'h90;
    assign sbox_data[151] = 8'h88;
    assign sbox_data[152] = 8'h46;
    assign sbox_data[153] = 8'hee;
    assign sbox_data[154] = 8'hb8;
    assign sbox_data[155] = 8'h14;
    assign sbox_data[156] = 8'hde;
    assign sbox_data[157] = 8'h5e;
    assign sbox_data[158] = 8'h0b;
    assign sbox_data[159] = 8'hdb;
    assign sbox_data[160] = 8'he0;
    assign sbox_data[161] = 8'h32;
    assign sbox_data[162] = 8'h3a;
    assign sbox_data[163] = 8'h0a;
    assign sbox_data[164] = 8'h49;
    assign sbox_data[165] = 8'h06;
    assign sbox_data[166] = 8'h24;
    assign sbox_data[167] = 8'h5c;
    assign sbox_data[168] = 8'hc2;
    assign sbox_data[169] = 8'hd3;
    assign sbox_data[170] = 8'hac;
    assign sbox_data[171] = 8'h62;
    assign sbox_data[172] = 8'h91;
    assign sbox_data[173] = 8'h95;
    assign sbox_data[174] = 8'he4;
    assign sbox_data[175] = 8'h79;
    assign sbox_data[176] = 8'he7;
    assign sbox_data[177] = 8'hc8;
    assign sbox_data[178] = 8'h37;
    assign sbox_data[179] = 8'h6d;
    assign sbox_data[180] = 8'h8d;
    assign sbox_data[181] = 8'hd5;
    assign sbox_data[182] = 8'h4e;
    assign sbox_data[183] = 8'ha9;
    assign sbox_data[184] = 8'h6c;
    assign sbox_data[185] = 8'h56;
    assign sbox_data[186] = 8'hf4;
    assign sbox_data[187] = 8'hea;
    assign sbox_data[188] = 8'h65;
    assign sbox_data[189] = 8'h7a;
    assign sbox_data[190] = 8'hae;
    assign sbox_data[191] = 8'h08;
    assign sbox_data[192] = 8'hba;
    assign sbox_data[193] = 8'h78;
    assign sbox_data[194] = 8'h25;
    assign sbox_data[195] = 8'h2e;
    assign sbox_data[196] = 8'h1c;
    assign sbox_data[197] = 8'ha6;
    assign sbox_data[198] = 8'hb4;
    assign sbox_data[199] = 8'hc6;
    assign sbox_data[200] = 8'he8;
    assign sbox_data[201] = 8'hdd;
    assign sbox_data[202] = 8'h74;
    assign sbox_data[203] = 8'h1f;
    assign sbox_data[204] = 8'h4b;
    assign sbox_data[205] = 8'hbd;
    assign sbox_data[206] = 8'h8b;
    assign sbox_data[207] = 8'h8a;
    assign sbox_data[208] = 8'h70;
    assign sbox_data[209] = 8'h3e;
    assign sbox_data[210] = 8'hb5;
    assign sbox_data[211] = 8'h66;
    assign sbox_data[212] = 8'h48;
    assign sbox_data[213] = 8'h03;
    assign sbox_data[214] = 8'hf6;
    assign sbox_data[215] = 8'h0e;
    assign sbox_data[216] = 8'h61;
    assign sbox_data[217] = 8'h35;
    assign sbox_data[218] = 8'h57;
    assign sbox_data[219] = 8'hb9;
    assign sbox_data[220] = 8'h86;
    assign sbox_data[221] = 8'hc1;
    assign sbox_data[222] = 8'h1d;
    assign sbox_data[223] = 8'h9e;
    assign sbox_data[224] = 8'he1;
    assign sbox_data[225] = 8'hf8;
    assign sbox_data[226] = 8'h98;
    assign sbox_data[227] = 8'h11;
    assign sbox_data[228] = 8'h69;
    assign sbox_data[229] = 8'hd9;
    assign sbox_data[230] = 8'h8e;
    assign sbox_data[231] = 8'h94;
    assign sbox_data[232] = 8'h9b;
    assign sbox_data[233] = 8'h1e;
    assign sbox_data[234] = 8'h87;
    assign sbox_data[235] = 8'he9;
    assign sbox_data[236] = 8'hce;
    assign sbox_data[237] = 8'h55;
    assign sbox_data[238] = 8'h28;
    assign sbox_data[239] = 8'hdf;
    assign sbox_data[240] = 8'h8c;
    assign sbox_data[241] = 8'ha1;
    assign sbox_data[242] = 8'h89;
    assign sbox_data[243] = 8'h0d;
    assign sbox_data[244] = 8'hbf;
    assign sbox_data[245] = 8'he6;
    assign sbox_data[246] = 8'h42;
    assign sbox_data[247] = 8'h68;
    assign sbox_data[248] = 8'h41;
    assign sbox_data[249] = 8'h99;
    assign sbox_data[250] = 8'h2d;
    assign sbox_data[251] = 8'h0f;
    assign sbox_data[252] = 8'hb0;
    assign sbox_data[253] = 8'h54;
    assign sbox_data[254] = 8'hbb;
    assign sbox_data[255] = 8'h16;
    
    // Output assignment
    assign out = sbox_data[index];

endmodule